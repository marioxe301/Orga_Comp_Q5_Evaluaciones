`define MIPS_AND 6'h24
`define MIPS_LW  6'h23
`define MIPS_BNE 6'h05